module AND_GATE
(
	input A,B,        // defining inputs A and B of AND gate 
	output C          // defining output of AND gate
);

assign C = A | B;   // Logic implementation
endmodule
